module main
(
input logic [1:0] button
)



endmodule